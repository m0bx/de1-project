library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity top_level is
    port (
         CLK   : in  std_logic;                       -- Main clock signal (e.g., 100 MHz)
         SW    : in  std_logic_vector(2 downto 0);   -- 16 physical switches (SW[1:0] determine mode, SW[2] determines if we are setting up the clock/alarm)
         CA    : out std_logic;                       -- active low
         CB    : out std_logic;                       
         CC    : out std_logic;                       
         CD    : out std_logic;                       
         CE    : out std_logic;                      
         CF    : out std_logic;                       
         CG    : out std_logic;                       
         DP    : out std_logic;                       -- Decimal point
         AN    : out std_logic_vector(7 downto 0);    -- 7-segment digit anode enables (active low)
         BTNC  : in  std_logic;                       -- stop/resume clock/alarm/stopwatch 
         BTND  : in  std_logic                        -- reset stopwatch
		 BTNL  : in  std_logic						  -- remove seconds/minutes from the counter (alarm or clock only)
		 BTNR  : in  std_logic						  -- add seconds/minutes from the counter (alarm or clock only)
    );
end entity top_level;

architecture behavioral of top_level is
    component bin2seg is
        port (
            clear : in  std_logic;
            bin   : in  std_logic_vector(3 downto 0);
            seg   : out std_logic_vector(6 downto 0)
        );
    end component;

    component display_mux is
        port (
             clk    : in  std_logic;
             rst    : in  std_logic;
             mode   : in  std_logic_vector(2 downto 0);
             digit0 : in  std_logic_vector(6 downto 0);
             digit1 : in  std_logic_vector(6 downto 0);
             digit2 : in  std_logic_vector(6 downto 0);
             digit3 : in  std_logic_vector(6 downto 0);
             digit4 : in  std_logic_vector(6 downto 0);
             digit5 : in  std_logic_vector(6 downto 0);
             digit6 : in  std_logic_vector(6 downto 0);
             digit7 : in  std_logic_vector(6 downto 0);
             -- seg    : out std_logic_vector(7 downto 0);  
             an     : out std_logic_vector(7 downto 0)
        );
    end component;

    signal disp_mode : std_logic_vector(2 downto 0);
    
    -- 4 bit binary value for each of the eight digits
    signal bin_digit0, bin_digit1, bin_digit2, bin_digit3,
           bin_digit4, bin_digit5, bin_digit6, bin_digit7 : std_logic_vector(3 downto 0);

    -- Seven-segment patterns generated by each bin2seg instance.
    signal sig_digit0, sig_digit1, sig_digit2, sig_digit3,
           sig_digit4, sig_digit5, sig_digit6, sig_digit7 : std_logic_vector(6 downto 0);

    -- multiplexer outputs 8-bit segment pattern and 8-bit anode enable.
    signal mux_seg : std_logic_vector(7 downto 0);
    signal mux_an  : std_logic_vector(7 downto 0);

begin

    disp_mode <= SW(2 downto 0);
    -- Digit value assignment.
    process(SW)
    begin
        case disp_mode is
            when "00"=>
                -- Clock only uses the first 4 digits. DP on 3rd AN is present
                bin_digit0 <= 
                bin_digit1 <= 
                bin_digit2 <= 
                bin_digit3 <= 
                -- Unused digits for Digital clock
                bin_digit4 <= "1111";
                bin_digit5 <= "1111";
                bin_digit6 <= "1111";
                bin_digit7 <= "1111";
              -- AN[2] will have DP enabled at all times
            when "10" =>
                -- stopwatch uses all 8 digits
                bin_digit0 <= 
                bin_digit1 <= 
                bin_digit2 <= 
                bin_digit3 <= 
                bin_digit4 <= 
                bin_digit5 <= 
                bin_digit6 <= 
                bin_digit7 <= 
				-- AN[4] will have DP enabled at all times (low active)
			when "01" =>
				-- Alarm
                bin_digit0 <= 
                bin_digit1 <= 
                bin_digit2 <= 
                bin_digit3 <= 
				-- Unused digits for alarm
                bin_digit4 <= "1111";
                bin_digit5 <= "1111";
                bin_digit6 <= "1111";
                bin_digit7 <= "1111";
            when others =>
                -- "11": Off mode. (Even though the display_mux blanks the output,
                -- you can assign any dummy value here.)
                bin_digit0 <= (others => '0');
                bin_digit1 <= (others => '0');
                bin_digit2 <= (others => '0');
                bin_digit3 <= (others => '0');
                bin_digit4 <= (others => '0');
                bin_digit5 <= (others => '0');
                bin_digit6 <= (others => '0');
                bin_digit7 <= (others => '0');
        end case;
    end process;

    u_display_mux: display_mux port map (
         clk    => CLK,        -- Scanning clock (should be divided from the system clock)
         rst    => BTNC,       -- Reset signal
         mode   => disp_mode,  -- Mode selection from SW(1 downto 0)
         digit0 => sig_digit0,
         digit1 => sig_digit1,
         digit2 => sig_digit2,
         digit3 => sig_digit3,
         digit4 => sig_digit4,
         digit5 => sig_digit5,
         digit6 => sig_digit6,
         digit7 => sig_digit7,
         seg    => mux_seg,    -- 8-bit segment output (MSB = DP)
         an     => mux_an      -- Anode (digit enable) outputs for each of the 8 digits
    );

-- mapping mux
    DP <= mux_seg(7);
    CA <= mux_seg(6);
    CB <= mux_seg(5);
    CC <= mux_seg(4);
    CD <= mux_seg(3);
    CE <= mux_seg(2);
    CF <= mux_seg(1);
    CG <= mux_seg(0);
    AN <= mux_an;

end architecture behavioral;
